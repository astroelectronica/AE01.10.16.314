.title KiCad schematic
.include "models/C2012X7R2A104K125AE_p.mod"
.include "models/INA188.lib"
XU2 /INP /INN VEE VDD VSS /GAIN1 /GAIN2 /OUT INA188
R4 /GAIN1 /GAIN2 12.4k
R2 /INN /INP 4.87k
R1 /IN /INN 100k
R3 /INP 0 20
V2 /IN 0 {VIN}
R5 /OUT 0 100k
V1 VDD 0 15
V3 0 VSS 15
V4 VEE 0 2.5
XU3 VSS 0 C2012X7R2A104K125AE_p
XU1 0 VDD C2012X7R2A104K125AE_p
XU4 0 VEE C2012X7R2A104K125AE_p
.end
